library verilog;
use verilog.vl_types.all;
entity alarma_vlg_vec_tst is
end alarma_vlg_vec_tst;
